package renacuajo_types;
    typedef logic[31:0] bus32_t;
    typedef logic[4:0] reg_addr_t;

    typedef logic[31:0] reg_t;

endpackage